module clk_div();

endmodule